/*
 * Created by 
   ../bin/Linux-x86_64-O/oasysGui 19.2-p002 on Fri Dec 24 14:38:39 2021
 * (C) Mentor Graphics Corporation
 */
/* CheckSum: 3486446019 */

module keep_H_C_value(clk, Rst, SFD, SRD, SW, SFA, ST, fdoor, rdoor, winbuzz, 
      alarmbuzz, heater, cooler, display);
   input clk;
   input Rst;
   input SFD;
   input SRD;
   input SW;
   input SFA;
   input [6:0]ST;
   output fdoor;
   output rdoor;
   output winbuzz;
   output alarmbuzz;
   output heater;
   output cooler;
   output [2:0]display;

   wire n_0_1_0;
   wire n_0_2_0;
   wire n_0_2_1;
   wire n_0_3_0;
   wire n_0_4_0;
   wire n_0_4_1;
   wire n_0_4_2;
   wire n_0_1;
   wire n_0_5_0;
   wire n_0_0;
   wire n_0_2;
   wire n_0_3;
   wire n_0_5_1;
   wire n_0_5_2;
   wire n_0_5_3;
   wire n_0_5_4;
   wire n_0_5_5;
   wire n_0_5_6;
   wire n_0_5_7;
   wire n_0_5_8;
   wire n_0_5_9;
   wire n_0_5_10;
   wire n_0_5_11;
   wire n_0_4;
   wire n_0_5_12;
   wire n_0_5_13;
   wire n_0_5_14;
   wire n_0_5_15;
   wire n_0_5_16;
   wire n_0_5_17;
   wire n_0_5_18;
   wire n_0_5_19;
   wire n_0_5;
   wire n_0_5_20;
   wire n_0_5_21;
   wire n_0_5_22;
   wire n_0_5_23;
   wire n_0_5_24;
   wire n_0_5_25;
   wire n_0_5_26;
   wire n_0_5_27;
   wire n_0_5_28;
   wire n_0_5_29;
   wire n_0_5_30;
   wire n_0_5_31;
   wire n_0_5_32;
   wire n_0_5_33;
   wire n_0_5_34;
   wire n_0_5_35;
   wire n_0_5_36;
   wire n_0_5_37;
   wire n_0_5_38;
   wire n_0_5_39;
   wire n_0_5_40;
   wire n_0_5_41;
   wire n_0_5_42;
   wire n_0_5_43;
   wire n_0_5_44;
   wire n_0_5_45;
   wire n_0_5_46;
   wire n_0_5_47;
   wire n_0_5_48;
   wire n_0_5_49;
   wire n_0_5_50;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;

   DFF_X2 \current_state_reg[1]  (.D(n_0_4), .CK(clk), .Q(display[1]), .QN());
   DFF_X2 \current_state_reg[2]  (.D(n_0_5), .CK(clk), .Q(display[2]), .QN());
   DFF_X2 \current_state_reg[0]  (.D(n_0_3), .CK(clk), .Q(display[0]), .QN());
   DLH_X1 cooler_reg (.D(n_0_2), .G(n_0_1), .Q(cooler));
   DLH_X1 heater_reg (.D(n_0_0), .G(n_0_1), .Q(heater));
   NAND2_X1 i_0_1_0 (.A1(display[1]), .A2(display[0]), .ZN(n_0_1_0));
   NOR2_X1 i_0_1_1 (.A1(n_0_1_0), .A2(display[2]), .ZN(alarmbuzz));
   NOR2_X1 i_0_2_0 (.A1(n_0_2_0), .A2(display[1]), .ZN(winbuzz));
   NAND2_X1 i_0_2_1 (.A1(display[2]), .A2(n_0_2_1), .ZN(n_0_2_0));
   INV_X1 i_0_2_2 (.A(display[0]), .ZN(n_0_2_1));
   INV_X1 i_0_3_0 (.A(display[1]), .ZN(n_0_3_0));
   NOR2_X1 i_0_3_1 (.A1(n_0_3_0), .A2(display[0]), .ZN(rdoor));
   INV_X1 i_0_4_0 (.A(n_0_4_0), .ZN(fdoor));
   NAND3_X1 i_0_4_1 (.A1(n_0_4_2), .A2(n_0_4_1), .A3(display[0]), .ZN(n_0_4_0));
   INV_X1 i_0_4_2 (.A(display[1]), .ZN(n_0_4_1));
   INV_X1 i_0_4_3 (.A(display[2]), .ZN(n_0_4_2));
   OAI21_X1 i_0_5_0 (.A(n_0_5_0), .B1(n_0_5_25), .B2(n_0_5_22), .ZN(n_0_1));
   NOR2_X1 i_0_5_1 (.A1(n_0_2), .A2(n_0_0), .ZN(n_0_5_0));
   NOR3_X1 i_0_5_2 (.A1(n_0_5_46), .A2(n_0_5_44), .A3(n_0_7), .ZN(n_0_0));
   NOR3_X1 i_0_5_3 (.A1(n_0_5_46), .A2(n_0_5_45), .A3(n_0_8), .ZN(n_0_2));
   NOR2_X1 i_0_5_4 (.A1(Rst), .A2(n_0_5_1), .ZN(n_0_3));
   AOI211_X1 i_0_5_5 (.A(n_0_5_8), .B(n_0_5_2), .C1(n_0_5_16), .C2(n_0_5_6), 
      .ZN(n_0_5_1));
   NOR3_X1 i_0_5_6 (.A1(n_0_6), .A2(n_0_5_4), .A3(n_0_5_3), .ZN(n_0_5_2));
   AOI21_X1 i_0_5_7 (.A(SFA), .B1(n_0_5_47), .B2(n_0_5_15), .ZN(n_0_5_3));
   AOI21_X1 i_0_5_8 (.A(n_0_5_5), .B1(n_0_7), .B2(n_0_5_44), .ZN(n_0_5_4));
   NOR3_X1 i_0_5_9 (.A1(n_0_7), .A2(n_0_5_44), .A3(SRD), .ZN(n_0_5_5));
   AOI21_X1 i_0_5_10 (.A(n_0_5_7), .B1(n_0_5_44), .B2(n_0_5_22), .ZN(n_0_5_6));
   AOI21_X1 i_0_5_11 (.A(n_0_5_41), .B1(n_0_5_28), .B2(n_0_5_11), .ZN(n_0_5_7));
   NOR3_X1 i_0_5_12 (.A1(n_0_5_34), .A2(n_0_5_9), .A3(n_0_5_18), .ZN(n_0_5_8));
   AOI21_X1 i_0_5_13 (.A(n_0_5_11), .B1(n_0_5_41), .B2(n_0_5_10), .ZN(n_0_5_9));
   NOR2_X1 i_0_5_14 (.A1(SRD), .A2(SW), .ZN(n_0_5_10));
   OAI21_X1 i_0_5_15 (.A(n_0_5_49), .B1(SRD), .B2(n_0_5_48), .ZN(n_0_5_11));
   NOR3_X1 i_0_5_16 (.A1(n_0_5_13), .A2(n_0_5_12), .A3(Rst), .ZN(n_0_4));
   NOR3_X1 i_0_5_17 (.A1(SRD), .A2(n_0_5_27), .A3(SFA), .ZN(n_0_5_12));
   AOI221_X1 i_0_5_18 (.A(n_0_5_17), .B1(n_0_5_39), .B2(n_0_5_37), .C1(n_0_5_16), 
      .C2(n_0_5_14), .ZN(n_0_5_13));
   INV_X1 i_0_5_19 (.A(n_0_5_15), .ZN(n_0_5_14));
   OAI21_X1 i_0_5_20 (.A(n_0_5_40), .B1(n_0_5_49), .B2(n_0_5_27), .ZN(n_0_5_15));
   OAI21_X1 i_0_5_21 (.A(n_0_5_22), .B1(SW), .B2(n_0_5_38), .ZN(n_0_5_16));
   AOI211_X1 i_0_5_22 (.A(n_0_5_33), .B(n_0_5_18), .C1(n_0_5_48), .C2(n_0_5_19), 
      .ZN(n_0_5_17));
   OAI21_X1 i_0_5_23 (.A(n_0_5_22), .B1(n_0_5_45), .B2(n_0_5_23), .ZN(n_0_5_18));
   AOI21_X1 i_0_5_24 (.A(SRD), .B1(n_0_5_47), .B2(n_0_5_40), .ZN(n_0_5_19));
   NOR3_X1 i_0_5_25 (.A1(n_0_5_24), .A2(n_0_5_20), .A3(Rst), .ZN(n_0_5));
   INV_X1 i_0_5_26 (.A(n_0_5_21), .ZN(n_0_5_20));
   OAI21_X1 i_0_5_27 (.A(n_0_5_31), .B1(n_0_5_26), .B2(n_0_5_22), .ZN(n_0_5_21));
   NAND2_X1 i_0_5_28 (.A1(n_0_5_45), .A2(n_0_5_23), .ZN(n_0_5_22));
   NOR2_X1 i_0_5_29 (.A1(n_0_5_46), .A2(n_0_8), .ZN(n_0_5_23));
   NOR3_X1 i_0_5_30 (.A1(SW), .A2(n_0_5_31), .A3(n_0_5_25), .ZN(n_0_5_24));
   INV_X1 i_0_5_31 (.A(n_0_5_26), .ZN(n_0_5_25));
   NOR2_X1 i_0_5_32 (.A1(n_0_5_41), .A2(n_0_5_27), .ZN(n_0_5_26));
   INV_X1 i_0_5_33 (.A(n_0_5_28), .ZN(n_0_5_27));
   OAI21_X1 i_0_5_34 (.A(ST[6]), .B1(n_0_5_30), .B2(n_0_5_29), .ZN(n_0_5_28));
   OR3_X1 i_0_5_35 (.A1(ST[4]), .A2(ST[3]), .A3(ST[5]), .ZN(n_0_5_29));
   AND3_X1 i_0_5_36 (.A1(ST[1]), .A2(ST[0]), .A3(ST[2]), .ZN(n_0_5_30));
   AOI22_X1 i_0_5_37 (.A1(n_0_5_39), .A2(n_0_5_36), .B1(n_0_5_48), .B2(n_0_5_32), 
      .ZN(n_0_5_31));
   NOR3_X1 i_0_5_38 (.A1(n_0_5_35), .A2(n_0_5_33), .A3(SRD), .ZN(n_0_5_32));
   NOR2_X1 i_0_5_39 (.A1(n_0_5_49), .A2(n_0_5_34), .ZN(n_0_5_33));
   NOR2_X1 i_0_5_40 (.A1(n_0_6), .A2(n_0_5_44), .ZN(n_0_5_34));
   NOR3_X1 i_0_5_41 (.A1(n_0_5_46), .A2(n_0_5_45), .A3(n_0_5_44), .ZN(n_0_5_35));
   INV_X1 i_0_5_42 (.A(n_0_5_37), .ZN(n_0_5_36));
   NOR2_X1 i_0_5_43 (.A1(n_0_5_48), .A2(n_0_8), .ZN(n_0_5_37));
   INV_X1 i_0_5_44 (.A(n_0_5_39), .ZN(n_0_5_38));
   NOR2_X1 i_0_5_45 (.A1(n_0_6), .A2(n_0_5_45), .ZN(n_0_5_39));
   INV_X1 i_0_5_46 (.A(n_0_5_41), .ZN(n_0_5_40));
   AOI21_X1 i_0_5_47 (.A(ST[6]), .B1(ST[5]), .B2(n_0_5_42), .ZN(n_0_5_41));
   NOR2_X1 i_0_5_48 (.A1(n_0_5_50), .A2(n_0_5_43), .ZN(n_0_5_42));
   NOR3_X1 i_0_5_49 (.A1(ST[2]), .A2(ST[1]), .A3(ST[3]), .ZN(n_0_5_43));
   INV_X1 i_0_5_50 (.A(n_0_8), .ZN(n_0_5_44));
   INV_X1 i_0_5_51 (.A(n_0_7), .ZN(n_0_5_45));
   INV_X1 i_0_5_52 (.A(n_0_6), .ZN(n_0_5_46));
   INV_X1 i_0_5_53 (.A(SW), .ZN(n_0_5_47));
   INV_X1 i_0_5_54 (.A(SFA), .ZN(n_0_5_48));
   INV_X1 i_0_5_55 (.A(SFD), .ZN(n_0_5_49));
   INV_X1 i_0_5_56 (.A(ST[4]), .ZN(n_0_5_50));
   BUF_X1 rt_shieldBuf__1 (.A(display[2]), .Z(n_0_6));
   BUF_X1 rt_shieldBuf__1__1__0 (.A(display[1]), .Z(n_0_7));
   BUF_X1 rt_shieldBuf__1__1__1 (.A(display[0]), .Z(n_0_8));
endmodule
