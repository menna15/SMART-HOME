/*
 * Created by 
   ../bin/Linux-x86_64-O/oasysGui 19.2-p002 on Fri Dec 24 14:52:53 2021
 * (C) Mentor Graphics Corporation
 */
/* CheckSum: 981913581 */

module Mealy(clk, Rst, SFD, SRD, SW, SFA, ST, fdoor, rdoor, winbuzz, alarmbuzz, 
      heater, cooler, display);
   input clk;
   input Rst;
   input SFD;
   input SRD;
   input SW;
   input SFA;
   input [6:0]ST;
   output fdoor;
   output rdoor;
   output winbuzz;
   output alarmbuzz;
   output heater;
   output cooler;
   output [2:0]display;

   wire [2:0]state;
   wire n_0_0_0;
   wire n_0_0_1;
   wire n_0_0_2;
   wire n_0_0;
   wire n_0_0_3;
   wire n_0_0_4;
   wire n_0_0_5;
   wire n_0_0_6;
   wire n_0_2_0;
   wire n_0_2_1;
   wire n_0_2_2;
   wire n_0_2_3;
   wire n_0_2_4;
   wire n_0_2_5;
   wire n_0_2_7;
   wire n_0_2_8;
   wire n_0_2_9;
   wire n_0_2_10;
   wire n_0_2_11;
   wire n_0_2_12;
   wire n_0_2_13;
   wire n_0_2_16;
   wire n_0_2_17;
   wire n_0_2_18;
   wire n_0_2_19;
   wire n_0_2_20;
   wire n_0_2_21;
   wire n_0_2_22;
   wire n_0_2_23;
   wire n_0_2_24;
   wire n_0_2_25;
   wire n_0_2_6;
   wire n_0_2_14;
   wire n_0_2_15;
   wire n_0_4_0;
   wire n_0_4_5;
   wire n_0_4_6;
   wire n_0_4_7;
   wire n_0_4_1;
   wire n_0_4_2;
   wire n_0_4_3;
   wire n_0_4_4;
   wire n_0_4_9;
   wire n_0_4_11;
   wire n_0_4_8;
   wire n_0_4_17;
   wire n_0_4_19;
   wire n_0_4_20;
   wire n_0_4_21;
   wire n_0_4_22;
   wire n_0_4_23;
   wire n_0_4_16;
   wire n_0_4_18;
   wire n_0_4_24;
   wire n_0_4_25;
   wire n_0_4_26;
   wire n_0_4_27;
   wire n_0_4_10;
   wire n_0_4_12;
   wire n_0_4_13;
   wire n_0_4_14;
   wire n_0_4_15;
   wire n_0_5_0;
   wire n_0_5_1;
   wire n_0_5_2;
   wire n_0_5_3;
   wire n_0_5_4;
   wire n_0_5_10;
   wire n_0_5_11;
   wire n_0_5_12;
   wire n_0_5_13;
   wire n_0_5_14;
   wire n_0_5_15;
   wire n_0_5_16;
   wire n_0_5_17;
   wire n_0_5_18;
   wire n_0_5_19;
   wire n_0_5_20;
   wire n_0_5_21;
   wire n_0_5_6;
   wire n_0_5_5;
   wire n_0_5_7;
   wire n_0_5_8;
   wire n_0_5_9;
   wire n_0_5_22;
   wire n_0_5_23;
   wire n_0_5_24;
   wire n_0_5_25;
   wire n_0_6_0;
   wire n_0_6_1;
   wire n_0_6_2;
   wire n_0_6_3;
   wire n_0_6_4;
   wire n_0_6_5;
   wire n_0_6_6;
   wire n_0_6_7;
   wire n_0_6_8;
   wire n_0_6_9;
   wire n_0_6_10;
   wire n_0_6_11;
   wire n_0_6_12;
   wire n_0_6_13;
   wire n_0_6_14;
   wire n_0_6_15;
   wire n_0_6_16;
   wire n_0_6_17;
   wire n_0_6_18;
   wire n_0_6_19;
   wire n_0_7_0;
   wire n_0_7_1;
   wire n_0_7_2;
   wire n_0_7_3;
   wire n_0_7_4;
   wire n_0_7_5;
   wire n_0_7_6;
   wire n_0_7_10;
   wire n_0_7_11;
   wire n_0_7_12;
   wire n_0_7_13;
   wire n_0_7_14;
   wire n_0_7_7;
   wire n_0_7_9;
   wire n_0_7_8;
   wire n_0_9_0;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_1_0;
   wire n_0_1_2;
   wire n_0_1_4;
   wire n_0_1_5;
   wire n_0_1_6;
   wire n_0_1_7;
   wire n_0_1_8;
   wire n_0_1_3;
   wire n_0_1_9;
   wire n_0_1_20;
   wire n_0_1_14;
   wire n_0_1_36;
   wire n_0_1_38;
   wire n_0_1_39;
   wire n_0_1_40;
   wire n_0_1_15;
   wire n_0_1_1;
   wire n_0_1_43;
   wire n_0_1_44;
   wire n_0_1_45;
   wire n_0_1_51;
   wire n_0_1_52;
   wire n_0_1_53;
   wire n_0_1_54;
   wire n_0_1_55;
   wire n_0_1_17;
   wire n_0_1_58;
   wire n_0_1_59;
   wire n_0_1_60;
   wire n_0_1_66;
   wire n_0_1_10;
   wire n_0_1_68;
   wire n_0_1_71;
   wire n_0_1_72;
   wire n_0_1_73;
   wire n_0_1_74;
   wire n_0_1_75;
   wire n_0_1_76;
   wire n_0_1_77;
   wire n_0_1_78;
   wire n_0_1_79;
   wire n_0_1_80;
   wire n_0_1_11;
   wire n_0_1_82;
   wire n_0_1_83;
   wire n_0_1_84;
   wire n_0_1_89;
   wire n_0_1_18;
   wire n_0_1_37;
   wire n_0_1_64;
   wire n_0_1_98;
   wire n_0_1_99;
   wire n_0_1_100;
   wire n_0_1_101;
   wire n_0_1_102;
   wire n_0_1_103;
   wire n_0_1_104;
   wire n_0_1_105;
   wire n_0_1_106;
   wire n_0_1_107;
   wire n_0_1_108;
   wire n_0_1_116;
   wire n_0_1_110;
   wire n_0_1_111;
   wire n_0_1_112;
   wire n_0_1_19;
   wire n_0_1_114;
   wire n_0_1_115;
   wire n_0_1;
   wire n_0_1_21;
   wire n_0_1_118;
   wire n_0_1_22;
   wire n_0_1_23;
   wire n_0_1_24;
   wire n_0_1_13;
   wire n_0_1_57;
   wire n_0_1_16;
   wire n_0_1_27;
   wire n_0_1_70;
   wire n_0_1_61;
   wire n_0_1_63;
   wire n_0_1_124;
   wire n_0_1_29;
   wire n_0_1_30;
   wire n_0_1_32;
   wire n_0_1_41;
   wire n_0_1_42;
   wire n_0_1_56;
   wire n_0_1_87;
   wire n_0_1_88;
   wire n_0_1_90;
   wire n_0_1_113;
   wire n_0_1_117;
   wire n_0_1_120;
   wire n_0_1_121;
   wire n_0_1_123;
   wire n_0_1_125;
   wire n_0_1_126;
   wire n_0_1_127;
   wire n_0_1_25;
   wire n_0_1_26;
   wire n_0_1_28;
   wire n_0_1_31;
   wire n_0_1_35;
   wire n_0_1_46;
   wire n_0_1_47;
   wire n_0_1_48;
   wire n_0_1_50;
   wire n_0_1_65;
   wire n_0_1_67;
   wire n_0_1_134;
   wire n_0_1_135;
   wire n_0_1_12;
   wire n_0_1_33;
   wire n_0_1_62;
   wire n_0_1_34;
   wire n_0_1_69;
   wire n_0_1_49;
   wire n_0_1_91;
   wire n_0_1_92;
   wire n_0_1_109;
   wire n_0_1_119;
   wire n_0_1_122;
   wire n_0_1_128;
   wire n_0_1_130;
   wire n_0_1_131;
   wire n_0_1_132;
   wire n_0_1_133;
   wire n_0_1_93;
   wire n_0_1_81;
   wire n_0_1_96;
   wire n_0_1_97;
   wire n_0_1_136;
   wire n_0_1_85;
   wire n_0_1_86;
   wire n_0_1_94;
   wire n_0_1_95;
   wire n_0_1_129;
   wire n_0_1_137;
   wire n_0_1_138;

   DFF_X2 \state_reg[0]  (.D(n_0_2), .CK(clk), .Q(state[0]), .QN());
   DFF_X2 \state_reg[2]  (.D(n_0_4), .CK(clk), .Q(state[2]), .QN());
   DFF_X2 \state_reg[1]  (.D(n_0_3), .CK(clk), .Q(state[1]), .QN());
   INV_X1 i_0_0_0 (.A(ST[1]), .ZN(n_0_0_0));
   INV_X1 i_0_0_1 (.A(ST[2]), .ZN(n_0_0_1));
   INV_X1 i_0_0_2 (.A(ST[3]), .ZN(n_0_0_2));
   INV_X1 i_0_0_3 (.A(n_0_0_3), .ZN(n_0_0));
   NAND2_X1 i_0_0_4 (.A1(n_0_0_4), .A2(n_0_0_6), .ZN(n_0_0_3));
   NAND3_X1 i_0_0_5 (.A1(n_0_0_5), .A2(ST[5]), .A3(ST[4]), .ZN(n_0_0_4));
   NAND3_X1 i_0_0_6 (.A1(n_0_0_1), .A2(n_0_0_0), .A3(n_0_0_2), .ZN(n_0_0_5));
   INV_X1 i_0_0_7 (.A(ST[6]), .ZN(n_0_0_6));
   INV_X1 i_0_2_0 (.A(n_0_0), .ZN(n_0_2_0));
   INV_X1 i_0_2_1 (.A(n_0_1), .ZN(n_0_2_1));
   INV_X1 i_0_2_2 (.A(SRD), .ZN(n_0_2_2));
   INV_X1 i_0_2_3 (.A(SFD), .ZN(n_0_2_3));
   NAND3_X1 i_0_2_4 (.A1(n_0_2_2), .A2(n_0_2_3), .A3(SFA), .ZN(n_0_2_4));
   INV_X1 i_0_2_5 (.A(n_0_2_4), .ZN(n_0_2_5));
   NAND2_X1 i_0_2_6 (.A1(n_0_2_5), .A2(n_0_2_6), .ZN(n_0_2_7));
   INV_X1 i_0_2_8 (.A(SW), .ZN(n_0_2_8));
   NAND4_X1 i_0_2_9 (.A1(n_0_2_8), .A2(n_0_2_2), .A3(n_0_2_3), .A4(SFA), 
      .ZN(n_0_2_9));
   OAI21_X1 i_0_2_7 (.A(n_0_2_7), .B1(state[2]), .B2(n_0_2_9), .ZN(n_0_2_10));
   INV_X1 i_0_2_10 (.A(state[2]), .ZN(n_0_2_11));
   INV_X1 i_0_2_11 (.A(state[1]), .ZN(n_0_2_12));
   NAND3_X1 i_0_2_13 (.A1(n_0_2_2), .A2(SFA), .A3(n_0_2_12), .ZN(n_0_2_13));
   NOR2_X1 i_0_2_12 (.A1(n_0_2_13), .A2(n_0_2_15), .ZN(n_0_2_16));
   NAND2_X1 i_0_2_14 (.A1(n_0_2_11), .A2(n_0_2_16), .ZN(n_0_2_17));
   NAND3_X1 i_0_2_19 (.A1(SFA), .A2(n_0_2_6), .A3(state[1]), .ZN(n_0_2_18));
   INV_X1 i_0_2_15 (.A(n_0_2_18), .ZN(n_0_2_19));
   NAND2_X1 i_0_2_16 (.A1(n_0_2_11), .A2(n_0_2_19), .ZN(n_0_2_20));
   XNOR2_X1 i_0_2_17 (.A(n_0_2_12), .B(state[0]), .ZN(n_0_2_21));
   NAND2_X1 i_0_2_18 (.A1(n_0_2_21), .A2(n_0_2_5), .ZN(n_0_2_22));
   NAND3_X1 i_0_2_20 (.A1(n_0_2_17), .A2(n_0_2_20), .A3(n_0_2_22), .ZN(n_0_2_23));
   NAND3_X1 i_0_2_21 (.A1(n_0_2_1), .A2(n_0_2_0), .A3(n_0_2_10), .ZN(n_0_2_24));
   INV_X1 i_0_2_22 (.A(n_0_2_23), .ZN(n_0_2_25));
   NAND2_X1 i_0_2_23 (.A1(n_0_2_24), .A2(n_0_2_25), .ZN(alarmbuzz));
   INV_X1 i_0_2_24 (.A(state[0]), .ZN(n_0_2_6));
   INV_X1 i_0_2_25 (.A(SFD), .ZN(n_0_2_14));
   NOR2_X1 i_0_2_26 (.A1(state[0]), .A2(n_0_2_14), .ZN(n_0_2_15));
   INV_X1 i_0_4_0 (.A(n_0_4_16), .ZN(n_0_4_0));
   INV_X1 i_0_4_11 (.A(SFD), .ZN(n_0_4_5));
   INV_X1 i_0_4_6 (.A(n_0_1), .ZN(n_0_4_6));
   INV_X1 i_0_4_8 (.A(n_0_0), .ZN(n_0_4_7));
   INV_X1 i_0_4_1 (.A(state[1]), .ZN(n_0_4_1));
   NAND2_X1 i_0_4_2 (.A1(n_0_4_1), .A2(n_0_4_4), .ZN(n_0_4_2));
   XNOR2_X1 i_0_4_3 (.A(state[1]), .B(state[0]), .ZN(n_0_4_3));
   INV_X1 i_0_4_9 (.A(state[2]), .ZN(n_0_4_4));
   NAND3_X1 i_0_4_7 (.A1(n_0_4_6), .A2(n_0_4_23), .A3(n_0_4_7), .ZN(n_0_4_9));
   NAND2_X1 i_0_4_18 (.A1(n_0_4_5), .A2(SRD), .ZN(n_0_4_11));
   INV_X1 i_0_4_20 (.A(n_0_4_11), .ZN(n_0_4_8));
   NAND2_X1 i_0_4_10 (.A1(n_0_4_9), .A2(n_0_4_15), .ZN(rdoor));
   NAND2_X1 i_0_4_4 (.A1(n_0_4_5), .A2(SRD), .ZN(n_0_4_17));
   INV_X1 i_0_4_5 (.A(SW), .ZN(n_0_4_19));
   NOR2_X1 i_0_4_13 (.A1(state[2]), .A2(n_0_4_19), .ZN(n_0_4_20));
   NOR2_X1 i_0_4_14 (.A1(n_0_4_17), .A2(n_0_4_20), .ZN(n_0_4_21));
   NAND2_X1 i_0_4_15 (.A1(n_0_4_27), .A2(n_0_4_21), .ZN(n_0_4_22));
   INV_X1 i_0_4_16 (.A(n_0_4_22), .ZN(n_0_4_23));
   NAND2_X1 i_0_4_12 (.A1(n_0_4_4), .A2(state[0]), .ZN(n_0_4_16));
   INV_X1 i_0_4_24 (.A(state[2]), .ZN(n_0_4_18));
   INV_X1 i_0_4_25 (.A(SFA), .ZN(n_0_4_24));
   NAND2_X1 i_0_4_17 (.A1(n_0_4_18), .A2(n_0_4_24), .ZN(n_0_4_25));
   NAND2_X1 i_0_4_19 (.A1(n_0_4_4), .A2(state[0]), .ZN(n_0_4_26));
   NAND3_X1 i_0_4_21 (.A1(n_0_4_25), .A2(n_0_4_26), .A3(state[1]), .ZN(n_0_4_27));
   NAND2_X1 i_0_4_22 (.A1(n_0_4_0), .A2(SRD), .ZN(n_0_4_10));
   INV_X1 i_0_4_23 (.A(n_0_4_8), .ZN(n_0_4_12));
   NAND2_X1 i_0_4_26 (.A1(n_0_4_10), .A2(n_0_4_12), .ZN(n_0_4_13));
   AOI22_X1 i_0_4_27 (.A1(n_0_4_3), .A2(n_0_4_2), .B1(n_0_4_2), .B2(n_0_4_4), 
      .ZN(n_0_4_14));
   NAND2_X1 i_0_4_28 (.A1(n_0_4_13), .A2(n_0_4_14), .ZN(n_0_4_15));
   INV_X1 i_0_5_0 (.A(n_0_0), .ZN(n_0_5_0));
   INV_X1 i_0_5_1 (.A(n_0_1), .ZN(n_0_5_1));
   INV_X1 i_0_5_2 (.A(SW), .ZN(n_0_5_2));
   OAI21_X1 i_0_5_3 (.A(SFD), .B1(n_0_5_2), .B2(state[2]), .ZN(n_0_5_3));
   INV_X1 i_0_5_4 (.A(state[2]), .ZN(n_0_5_4));
   NAND3_X1 i_0_5_5 (.A1(state[1]), .A2(state[0]), .A3(n_0_5_4), .ZN(n_0_5_10));
   AOI21_X1 i_0_5_6 (.A(n_0_5_3), .B1(n_0_5_25), .B2(n_0_5_10), .ZN(n_0_5_11));
   INV_X1 i_0_5_13 (.A(state[0]), .ZN(n_0_5_12));
   INV_X1 i_0_5_7 (.A(state[1]), .ZN(n_0_5_13));
   NAND3_X1 i_0_5_8 (.A1(SFD), .A2(n_0_5_13), .A3(state[2]), .ZN(n_0_5_14));
   NAND2_X1 i_0_5_9 (.A1(n_0_5_6), .A2(SFD), .ZN(n_0_5_15));
   NAND3_X1 i_0_5_10 (.A1(n_0_5_1), .A2(n_0_5_0), .A3(n_0_5_11), .ZN(n_0_5_16));
   NOR2_X1 i_0_5_11 (.A1(n_0_5_14), .A2(n_0_5_12), .ZN(n_0_5_17));
   INV_X1 i_0_5_12 (.A(n_0_5_15), .ZN(n_0_5_18));
   INV_X1 i_0_5_14 (.A(n_0_5_12), .ZN(n_0_5_19));
   NAND2_X1 i_0_5_15 (.A1(n_0_5_14), .A2(n_0_5_19), .ZN(n_0_5_20));
   AOI21_X1 i_0_5_16 (.A(n_0_5_17), .B1(n_0_5_18), .B2(n_0_5_20), .ZN(n_0_5_21));
   NAND2_X1 i_0_5_17 (.A1(n_0_5_16), .A2(n_0_5_21), .ZN(fdoor));
   XNOR2_X1 i_0_5_21 (.A(state[1]), .B(state[2]), .ZN(n_0_5_6));
   INV_X1 i_0_5_18 (.A(state[1]), .ZN(n_0_5_5));
   INV_X1 i_0_5_19 (.A(n_0_5_5), .ZN(n_0_5_7));
   NAND2_X1 i_0_5_20 (.A1(n_0_5_7), .A2(state[2]), .ZN(n_0_5_8));
   INV_X1 i_0_5_22 (.A(SRD), .ZN(n_0_5_9));
   NOR2_X1 i_0_5_23 (.A1(state[2]), .A2(n_0_5_9), .ZN(n_0_5_22));
   NAND2_X1 i_0_5_24 (.A1(n_0_5_5), .A2(n_0_5_22), .ZN(n_0_5_23));
   NAND2_X1 i_0_5_25 (.A1(n_0_5_4), .A2(SFA), .ZN(n_0_5_24));
   NAND3_X1 i_0_5_26 (.A1(n_0_5_8), .A2(n_0_5_23), .A3(n_0_5_24), .ZN(n_0_5_25));
   AOI21_X1 i_0_6_0 (.A(n_0_6_0), .B1(n_0_6_2), .B2(n_0_6_11), .ZN(cooler));
   NAND2_X1 i_0_6_1 (.A1(n_0_6_1), .A2(n_0_1), .ZN(n_0_6_0));
   INV_X1 i_0_6_2 (.A(n_0_0), .ZN(n_0_6_1));
   AOI21_X1 i_0_6_3 (.A(n_0_6_3), .B1(n_0_6_5), .B2(n_0_6_10), .ZN(n_0_6_2));
   INV_X1 i_0_6_4 (.A(n_0_6_4), .ZN(n_0_6_3));
   NAND3_X1 i_0_6_5 (.A1(n_0_6_19), .A2(n_0_6_17), .A3(state[2]), .ZN(n_0_6_4));
   INV_X1 i_0_6_6 (.A(n_0_6_6), .ZN(n_0_6_5));
   NAND4_X1 i_0_6_7 (.A1(n_0_6_9), .A2(n_0_6_8), .A3(n_0_6_7), .A4(n_0_6_15), 
      .ZN(n_0_6_6));
   INV_X1 i_0_6_8 (.A(SFD), .ZN(n_0_6_7));
   INV_X1 i_0_6_9 (.A(SRD), .ZN(n_0_6_8));
   INV_X1 i_0_6_10 (.A(SFA), .ZN(n_0_6_9));
   NAND2_X1 i_0_6_11 (.A1(state[1]), .A2(state[0]), .ZN(n_0_6_10));
   NAND3_X1 i_0_6_12 (.A1(n_0_6_18), .A2(n_0_6_16), .A3(n_0_6_12), .ZN(n_0_6_11));
   INV_X1 i_0_6_13 (.A(n_0_6_13), .ZN(n_0_6_12));
   NAND2_X1 i_0_6_14 (.A1(n_0_6_15), .A2(n_0_6_14), .ZN(n_0_6_13));
   INV_X1 i_0_6_15 (.A(state[2]), .ZN(n_0_6_14));
   INV_X1 i_0_6_16 (.A(SW), .ZN(n_0_6_15));
   OAI21_X1 i_0_6_17 (.A(n_0_6_17), .B1(n_0_6_19), .B2(SFA), .ZN(n_0_6_16));
   INV_X1 i_0_6_18 (.A(state[0]), .ZN(n_0_6_17));
   OAI21_X1 i_0_6_19 (.A(n_0_6_19), .B1(SFA), .B2(SRD), .ZN(n_0_6_18));
   INV_X1 i_0_6_20 (.A(state[1]), .ZN(n_0_6_19));
   INV_X1 i_0_7_0 (.A(n_0_7_0), .ZN(heater));
   NAND2_X1 i_0_7_1 (.A1(n_0_0), .A2(n_0_7_1), .ZN(n_0_7_0));
   OAI21_X1 i_0_7_2 (.A(n_0_7_2), .B1(n_0_7_6), .B2(n_0_7_3), .ZN(n_0_7_1));
   NAND3_X1 i_0_7_3 (.A1(n_0_7_12), .A2(n_0_7_11), .A3(state[2]), .ZN(n_0_7_2));
   OAI21_X1 i_0_7_4 (.A(n_0_7_5), .B1(n_0_7_4), .B2(n_0_7_7), .ZN(n_0_7_3));
   INV_X1 i_0_7_5 (.A(SFA), .ZN(n_0_7_4));
   INV_X1 i_0_7_6 (.A(SW), .ZN(n_0_7_5));
   AOI22_X1 i_0_7_7 (.A1(n_0_7_10), .A2(n_0_7_13), .B1(n_0_7_8), .B2(n_0_7_14), 
      .ZN(n_0_7_6));
   OAI21_X1 i_0_7_8 (.A(n_0_7_12), .B1(SRD), .B2(n_0_7_11), .ZN(n_0_7_10));
   INV_X1 i_0_7_9 (.A(state[0]), .ZN(n_0_7_11));
   INV_X1 i_0_7_10 (.A(state[1]), .ZN(n_0_7_12));
   INV_X1 i_0_7_11 (.A(state[2]), .ZN(n_0_7_13));
   INV_X1 i_0_7_15 (.A(SFD), .ZN(n_0_7_14));
   INV_X1 i_0_7_12 (.A(n_0_7_9), .ZN(n_0_7_7));
   NAND2_X1 i_0_7_13 (.A1(state[1]), .A2(state[0]), .ZN(n_0_7_9));
   AOI21_X1 i_0_7_14 (.A(SRD), .B1(state[1]), .B2(state[0]), .ZN(n_0_7_8));
   INV_X1 i_0_9_0 (.A(Rst), .ZN(n_0_9_0));
   AND2_X1 i_0_9_1 (.A1(n_0_9_0), .A2(display[0]), .ZN(n_0_2));
   AND2_X1 i_0_9_2 (.A1(n_0_9_0), .A2(display[1]), .ZN(n_0_3));
   AND2_X1 i_0_9_3 (.A1(n_0_9_0), .A2(display[2]), .ZN(n_0_4));
   INV_X1 i_0_1_0 (.A(n_0_0), .ZN(n_0_1_0));
   INV_X1 i_0_1_2 (.A(SFD), .ZN(n_0_1_2));
   NAND3_X1 i_0_1_1 (.A1(n_0_1_2), .A2(SW), .A3(n_0_1_22), .ZN(n_0_1_4));
   INV_X1 i_0_1_5 (.A(SFA), .ZN(n_0_1_5));
   INV_X1 i_0_1_6 (.A(SRD), .ZN(n_0_1_6));
   NAND2_X1 i_0_1_7 (.A1(n_0_1_5), .A2(n_0_1_6), .ZN(n_0_1_7));
   NOR2_X1 i_0_1_3 (.A1(n_0_1_4), .A2(n_0_1_7), .ZN(n_0_1_8));
   NAND2_X1 i_0_1_9 (.A1(SFD), .A2(state[2]), .ZN(n_0_1_3));
   INV_X1 i_0_1_18 (.A(state[1]), .ZN(n_0_1_9));
   NAND3_X1 i_0_1_4 (.A1(n_0_1_116), .A2(n_0_1_0), .A3(n_0_1_8), .ZN(n_0_1_20));
   NAND2_X1 i_0_1_8 (.A1(n_0_1_131), .A2(n_0_1_20), .ZN(winbuzz));
   XNOR2_X1 i_0_1_22 (.A(SFD), .B(n_0_1_35), .ZN(n_0_1_14));
   INV_X1 i_0_1_37 (.A(SFD), .ZN(n_0_1_36));
   NAND3_X1 i_0_1_19 (.A1(n_0_1_36), .A2(state[2]), .A3(n_0_1_22), .ZN(n_0_1_38));
   NAND3_X1 i_0_1_40 (.A1(SFD), .A2(n_0_1_22), .A3(n_0_1_35), .ZN(n_0_1_39));
   NAND2_X1 i_0_1_23 (.A1(n_0_1_38), .A2(n_0_1_39), .ZN(n_0_1_40));
   INV_X1 i_0_1_24 (.A(n_0_1_40), .ZN(n_0_1_15));
   NOR2_X1 i_0_1_44 (.A1(SFA), .A2(state[2]), .ZN(n_0_1_1));
   AOI21_X1 i_0_1_11 (.A(n_0_1_76), .B1(n_0_1_71), .B2(n_0_1_112), .ZN(
      display[0]));
   NAND3_X1 i_0_1_46 (.A1(n_0_1_44), .A2(n_0_1_69), .A3(state[1]), .ZN(n_0_1_43));
   NAND2_X1 i_0_1_47 (.A1(n_0_1_94), .A2(SW), .ZN(n_0_1_44));
   OAI21_X1 i_0_1_48 (.A(n_0_1_66), .B1(n_0_1_60), .B2(SFA), .ZN(n_0_1_45));
   NAND3_X1 i_0_1_12 (.A1(n_0_1_53), .A2(n_0_1_100), .A3(n_0_1_52), .ZN(n_0_1_51));
   NAND2_X1 i_0_1_55 (.A1(SFD), .A2(state[2]), .ZN(n_0_1_52));
   OAI21_X1 i_0_1_13 (.A(n_0_1_118), .B1(SFD), .B2(state[2]), .ZN(n_0_1_53));
   AOI21_X1 i_0_1_14 (.A(n_0_1_17), .B1(n_0_1_55), .B2(n_0_1_93), .ZN(n_0_1_54));
   INV_X1 i_0_1_15 (.A(n_0_1_1), .ZN(n_0_1_55));
   INV_X1 i_0_1_16 (.A(state[1]), .ZN(n_0_1_17));
   AOI21_X1 i_0_1_17 (.A(n_0_1_80), .B1(n_0_1_71), .B2(n_0_1_58), .ZN(display[2]));
   NOR2_X1 i_0_1_27 (.A1(n_0_1), .A2(n_0_1_59), .ZN(n_0_1_58));
   AOI21_X1 i_0_1_31 (.A(n_0_1_60), .B1(n_0_1_115), .B2(n_0_1_118), .ZN(n_0_1_59));
   INV_X1 i_0_1_43 (.A(SW), .ZN(n_0_1_60));
   INV_X1 i_0_1_70 (.A(SRD), .ZN(n_0_1_66));
   INV_X1 i_0_1_71 (.A(SFA), .ZN(n_0_1_10));
   AOI22_X1 i_0_1_45 (.A1(n_0_1_19), .A2(n_0_1_28), .B1(n_0_1_69), .B2(state[0]), 
      .ZN(n_0_1_68));
   INV_X1 i_0_1_52 (.A(n_0_0), .ZN(n_0_1_71));
   NAND2_X1 i_0_1_76 (.A1(n_0_1_19), .A2(n_0_1_10), .ZN(n_0_1_72));
   INV_X1 i_0_1_77 (.A(n_0_1_72), .ZN(n_0_1_73));
   NAND2_X1 i_0_1_21 (.A1(n_0_1_43), .A2(n_0_1_53), .ZN(n_0_1_74));
   INV_X1 i_0_1_29 (.A(n_0_1_47), .ZN(n_0_1_75));
   AOI21_X1 i_0_1_34 (.A(n_0_1_74), .B1(n_0_1_99), .B2(n_0_1_75), .ZN(n_0_1_76));
   INV_X1 i_0_1_56 (.A(n_0_1_86), .ZN(n_0_1_77));
   NAND2_X1 i_0_1_58 (.A1(n_0_1_100), .A2(n_0_1_46), .ZN(n_0_1_78));
   NAND2_X1 i_0_1_63 (.A1(n_0_1_68), .A2(n_0_1_46), .ZN(n_0_1_79));
   AOI21_X1 i_0_1_72 (.A(n_0_1_77), .B1(n_0_1_78), .B2(n_0_1_79), .ZN(n_0_1_80));
   NAND3_X1 i_0_1_85 (.A1(n_0_1_82), .A2(n_0_1_83), .A3(n_0_1_84), .ZN(n_0_1_11));
   NOR2_X1 i_0_1_86 (.A1(ST[5]), .A2(ST[3]), .ZN(n_0_1_82));
   NAND3_X1 i_0_1_87 (.A1(ST[1]), .A2(ST[2]), .A3(ST[0]), .ZN(n_0_1_83));
   INV_X1 i_0_1_88 (.A(ST[4]), .ZN(n_0_1_84));
   INV_X1 i_0_1_93 (.A(ST[6]), .ZN(n_0_1_89));
   NOR2_X1 i_0_1_94 (.A1(n_0_1_89), .A2(SW), .ZN(n_0_1_18));
   INV_X1 i_0_1_97 (.A(SFD), .ZN(n_0_1_37));
   INV_X1 i_0_1_99 (.A(n_0_1_60), .ZN(n_0_1_64));
   AOI22_X1 i_0_1_53 (.A1(n_0_1_125), .A2(n_0_1_101), .B1(n_0_1_100), .B2(
      n_0_1_136), .ZN(n_0_1_98));
   NAND2_X1 i_0_1_35 (.A1(n_0_1_45), .A2(n_0_1_52), .ZN(n_0_1_99));
   NAND2_X1 i_0_1_81 (.A1(n_0_1_10), .A2(n_0_1_66), .ZN(n_0_1_100));
   NAND3_X1 i_0_1_105 (.A1(n_0_1_102), .A2(n_0_1_103), .A3(n_0_1_104), .ZN(
      n_0_1_101));
   NOR2_X1 i_0_1_106 (.A1(ST[4]), .A2(ST[5]), .ZN(n_0_1_102));
   NAND3_X1 i_0_1_107 (.A1(ST[1]), .A2(ST[0]), .A3(ST[2]), .ZN(n_0_1_103));
   INV_X1 i_0_1_108 (.A(ST[3]), .ZN(n_0_1_104));
   NOR2_X1 i_0_1_109 (.A1(ST[4]), .A2(ST[5]), .ZN(n_0_1_105));
   NAND3_X1 i_0_1_110 (.A1(ST[1]), .A2(ST[0]), .A3(ST[2]), .ZN(n_0_1_106));
   INV_X1 i_0_1_111 (.A(ST[3]), .ZN(n_0_1_107));
   NAND3_X1 i_0_1_112 (.A1(n_0_1_105), .A2(n_0_1_106), .A3(n_0_1_107), .ZN(
      n_0_1_108));
   NAND2_X1 i_0_1_84 (.A1(n_0_1_108), .A2(ST[6]), .ZN(n_0_1_116));
   OAI22_X1 i_0_1_54 (.A1(n_0_1_98), .A2(n_0_0), .B1(n_0_1_54), .B2(n_0_1_51), 
      .ZN(display[1]));
   NAND2_X1 i_0_1_41 (.A1(n_0_1_42), .A2(n_0_1_19), .ZN(n_0_1_110));
   INV_X1 i_0_1_118 (.A(n_0_1_73), .ZN(n_0_1_111));
   NAND3_X1 i_0_1_50 (.A1(n_0_1_12), .A2(n_0_1_110), .A3(n_0_1_111), .ZN(
      n_0_1_112));
   INV_X1 i_0_1_120 (.A(SFD), .ZN(n_0_1_19));
   INV_X1 i_0_1_121 (.A(SFD), .ZN(n_0_1_114));
   NAND3_X1 i_0_1_104 (.A1(n_0_1_10), .A2(n_0_1_66), .A3(n_0_1_114), .ZN(
      n_0_1_115));
   INV_X1 i_0_1_113 (.A(n_0_1_116), .ZN(n_0_1));
   INV_X1 i_0_1_60 (.A(ST[6]), .ZN(n_0_1_21));
   NOR2_X1 i_0_1_61 (.A1(state[1]), .A2(state[0]), .ZN(n_0_1_118));
   INV_X1 i_0_1_32 (.A(state[0]), .ZN(n_0_1_22));
   INV_X1 i_0_1_26 (.A(state[2]), .ZN(n_0_1_23));
   NAND2_X1 i_0_1_10 (.A1(n_0_1_23), .A2(state[1]), .ZN(n_0_1_24));
   NAND2_X1 i_0_1_28 (.A1(n_0_1_23), .A2(state[1]), .ZN(n_0_1_13));
   NAND2_X1 i_0_1_96 (.A1(n_0_1_5), .A2(SW), .ZN(n_0_1_57));
   INV_X1 i_0_1_98 (.A(n_0_1_57), .ZN(n_0_1_16));
   NAND2_X1 i_0_1_30 (.A1(n_0_1_33), .A2(SRD), .ZN(n_0_1_27));
   INV_X1 i_0_1_101 (.A(SW), .ZN(n_0_1_70));
   NOR2_X1 i_0_1_33 (.A1(n_0_1_22), .A2(n_0_1_70), .ZN(n_0_1_61));
   INV_X1 i_0_1_25 (.A(n_0_1_24), .ZN(n_0_1_63));
   NAND2_X1 i_0_1_36 (.A1(n_0_1_22), .A2(state[1]), .ZN(n_0_1_124));
   INV_X1 i_0_1_38 (.A(n_0_1_124), .ZN(n_0_1_29));
   INV_X1 i_0_1_130 (.A(SRD), .ZN(n_0_1_30));
   INV_X1 i_0_1_57 (.A(n_0_1_17), .ZN(n_0_1_32));
   INV_X1 i_0_1_79 (.A(state[0]), .ZN(n_0_1_41));
   AOI21_X1 i_0_1_78 (.A(n_0_1_30), .B1(n_0_1_32), .B2(n_0_1_41), .ZN(n_0_1_42));
   NAND2_X1 i_0_1_73 (.A1(state[1]), .A2(state[0]), .ZN(n_0_1_56));
   NAND3_X1 i_0_1_74 (.A1(n_0_1_18), .A2(n_0_1_19), .A3(n_0_1_56), .ZN(n_0_1_87));
   NOR2_X1 i_0_1_90 (.A1(state[2]), .A2(SW), .ZN(n_0_1_88));
   INV_X1 i_0_1_91 (.A(state[1]), .ZN(n_0_1_90));
   INV_X1 i_0_1_92 (.A(state[0]), .ZN(n_0_1_113));
   NAND2_X1 i_0_1_122 (.A1(n_0_1_90), .A2(n_0_1_113), .ZN(n_0_1_117));
   INV_X1 i_0_1_124 (.A(n_0_1_21), .ZN(n_0_1_120));
   NAND3_X1 i_0_1_134 (.A1(n_0_1_88), .A2(n_0_1_117), .A3(n_0_1_120), .ZN(
      n_0_1_121));
   NAND3_X1 i_0_1_135 (.A1(n_0_1_48), .A2(n_0_1_120), .A3(state[2]), .ZN(
      n_0_1_123));
   NAND3_X1 i_0_1_59 (.A1(n_0_1_87), .A2(n_0_1_121), .A3(n_0_1_123), .ZN(
      n_0_1_125));
   NAND2_X1 i_0_1_39 (.A1(n_0_1_3), .A2(n_0_1_9), .ZN(n_0_1_126));
   INV_X1 i_0_1_42 (.A(n_0_1_126), .ZN(n_0_1_127));
   NAND2_X1 i_0_1_49 (.A1(n_0_1_15), .A2(n_0_1_127), .ZN(n_0_1_25));
   NAND2_X1 i_0_1_51 (.A1(n_0_1_14), .A2(n_0_1_29), .ZN(n_0_1_26));
   NAND2_X1 i_0_1_62 (.A1(state[1]), .A2(state[0]), .ZN(n_0_1_28));
   NAND2_X1 i_0_1_102 (.A1(state[1]), .A2(state[0]), .ZN(n_0_1_31));
   INV_X1 i_0_1_95 (.A(state[2]), .ZN(n_0_1_35));
   NAND2_X1 i_0_1_64 (.A1(n_0_1_48), .A2(state[2]), .ZN(n_0_1_46));
   INV_X1 i_0_1_20 (.A(n_0_1_31), .ZN(n_0_1_47));
   NOR2_X1 i_0_1_67 (.A1(state[1]), .A2(state[0]), .ZN(n_0_1_48));
   NOR2_X1 i_0_1_123 (.A1(n_0_1_10), .A2(state[2]), .ZN(n_0_1_50));
   NAND2_X1 i_0_1_115 (.A1(n_0_1_33), .A2(SRD), .ZN(n_0_1_65));
   NOR2_X1 i_0_1_119 (.A1(n_0_1_13), .A2(SFA), .ZN(n_0_1_67));
   INV_X1 i_0_1_133 (.A(ST[6]), .ZN(n_0_1_134));
   AOI21_X1 i_0_1_131 (.A(n_0_1_134), .B1(n_0_1_50), .B2(n_0_1_31), .ZN(
      n_0_1_135));
   NAND3_X1 i_0_1_132 (.A1(n_0_1_133), .A2(n_0_1_11), .A3(n_0_1_135), .ZN(
      n_0_1_12));
   NAND2_X1 i_0_1_128 (.A1(n_0_1_62), .A2(state[1]), .ZN(n_0_1_33));
   INV_X1 i_0_1_129 (.A(state[2]), .ZN(n_0_1_62));
   INV_X1 i_0_1_139 (.A(state[1]), .ZN(n_0_1_34));
   INV_X1 i_0_1_68 (.A(state[2]), .ZN(n_0_1_69));
   INV_X1 i_0_1_65 (.A(state[2]), .ZN(n_0_1_49));
   NAND3_X1 i_0_1_66 (.A1(n_0_1_49), .A2(state[1]), .A3(state[0]), .ZN(n_0_1_91));
   OAI21_X1 i_0_1_89 (.A(n_0_1_91), .B1(n_0_1_13), .B2(SFA), .ZN(n_0_1_92));
   NAND2_X1 i_0_1_125 (.A1(state[1]), .A2(state[0]), .ZN(n_0_1_109));
   NAND3_X1 i_0_1_126 (.A1(n_0_1_109), .A2(n_0_1_34), .A3(SRD), .ZN(n_0_1_119));
   NAND2_X1 i_0_1_144 (.A1(state[2]), .A2(SRD), .ZN(n_0_1_122));
   NAND3_X1 i_0_1_145 (.A1(n_0_1_92), .A2(n_0_1_119), .A3(n_0_1_122), .ZN(
      n_0_1_128));
   NAND3_X1 i_0_1_100 (.A1(n_0_1_25), .A2(n_0_1_128), .A3(n_0_1_26), .ZN(
      n_0_1_130));
   NAND2_X1 i_0_1_136 (.A1(n_0_1_138), .A2(n_0_1_130), .ZN(n_0_1_131));
   NOR2_X1 i_0_1_103 (.A1(state[1]), .A2(state[0]), .ZN(n_0_1_132));
   XNOR2_X1 i_0_1_116 (.A(n_0_1_132), .B(state[2]), .ZN(n_0_1_133));
   INV_X1 i_0_1_69 (.A(state[0]), .ZN(n_0_1_93));
   INV_X1 i_0_1_75 (.A(state[0]), .ZN(n_0_1_81));
   NAND2_X1 i_0_1_83 (.A1(n_0_1_17), .A2(n_0_1_37), .ZN(n_0_1_96));
   NAND2_X1 i_0_1_117 (.A1(n_0_1_69), .A2(n_0_1_37), .ZN(n_0_1_97));
   OAI21_X1 i_0_1_127 (.A(n_0_1_96), .B1(n_0_1_97), .B2(n_0_1_64), .ZN(n_0_1_136));
   NAND2_X1 i_0_1_80 (.A1(n_0_1_81), .A2(SFA), .ZN(n_0_1_85));
   NAND3_X1 i_0_1_114 (.A1(n_0_1_85), .A2(n_0_1_69), .A3(state[1]), .ZN(n_0_1_86));
   NAND2_X1 i_0_1_82 (.A1(n_0_1_81), .A2(SFA), .ZN(n_0_1_94));
   NAND3_X1 i_0_1_137 (.A1(n_0_1_67), .A2(n_0_1_65), .A3(SW), .ZN(n_0_1_95));
   NAND2_X1 i_0_1_138 (.A1(n_0_1_63), .A2(n_0_1_61), .ZN(n_0_1_129));
   NAND2_X1 i_0_1_140 (.A1(n_0_1_16), .A2(n_0_1_27), .ZN(n_0_1_137));
   NAND3_X1 i_0_1_141 (.A1(n_0_1_95), .A2(n_0_1_129), .A3(n_0_1_137), .ZN(
      n_0_1_138));
endmodule
