/*
 * Created by 
   ../bin/Linux-x86_64-O/oasysGui 19.2-p002 on Thu Dec 23 21:13:15 2021
 * (C) Mentor Graphics Corporation
 */
/* CheckSum: 607411740 */

module Mealy(clk, Rst, SFD, SRD, SW, SFA, ST, fdoor, rdoor, winbuzz, alarmbuzz, 
      heater, cooler, display);
   input clk;
   input Rst;
   input SFD;
   input SRD;
   input SW;
   input SFA;
   input [6:0]ST;
   output fdoor;
   output rdoor;
   output winbuzz;
   output alarmbuzz;
   output heater;
   output cooler;
   output [2:0]display;

   wire n_0_0_0;
   wire n_0_0_1;
   wire n_0_0_2;
   wire n_0_0;
   wire n_0_0_3;
   wire n_0_0_4;
   wire n_0_0_5;
   wire n_0_0_6;
   wire n_0_1_0;
   wire n_0_1_1;
   wire n_0_1_2;
   wire n_0_1_3;
   wire n_0_1_4;
   wire n_0_1_5;
   wire n_0_1_6;
   wire n_0_1_7;
   wire n_0_1_8;
   wire n_0_1_9;
   wire n_0_1_10;
   wire n_0_1_11;
   wire n_0_1_12;
   wire n_0_1_13;
   wire n_0_1_14;
   wire n_0_1_15;
   wire n_0_1_16;
   wire n_0_1_17;
   wire n_0_2_0;
   wire n_0_2_1;
   wire n_0_2_2;
   wire n_0_2_3;
   wire n_0_2_4;
   wire n_0_2_5;
   wire n_0_2_6;
   wire n_0_2_7;
   wire n_0_2_8;
   wire n_0_2_9;
   wire n_0_2_10;
   wire n_0_2_11;
   wire n_0_2_12;
   wire n_0_2_13;
   wire n_0_2_14;
   wire n_0_2_15;
   wire n_0_2_16;
   wire n_0_2_17;
   wire n_0_3_0;
   wire n_0_3_1;
   wire n_0_3_2;
   wire n_0_3_3;
   wire n_0_3_4;
   wire n_0_3_5;
   wire n_0_3_6;
   wire n_0_3_9;
   wire n_0_3_7;
   wire n_0_3_11;
   wire n_0_3_8;
   wire n_0_3_10;
   wire n_0_3_12;
   wire n_0_3_13;
   wire n_0_3_14;
   wire n_0_3_15;
   wire n_0_3_16;
   wire n_0_4_1;
   wire n_0_4_7;
   wire n_0_4_9;
   wire n_0_4_0;
   wire n_0_4_2;
   wire n_0_4_3;
   wire n_0_4_4;
   wire n_0_4_5;
   wire n_0_4_6;
   wire n_0_4_8;
   wire n_0_4_10;
   wire n_0_4_11;
   wire n_0_4_12;
   wire n_0_4_13;
   wire n_0_4_14;
   wire n_0_4_15;
   wire n_0_4_16;
   wire n_0_6_8;
   wire n_0_6_9;
   wire n_0_6_10;
   wire n_0_6_11;
   wire n_0_6_12;
   wire n_0_6_0;
   wire n_0_6_1;
   wire n_0_6_2;
   wire n_0_6_3;
   wire n_0_6_4;
   wire n_0_6_5;
   wire n_0_6_6;
   wire n_0_6_7;
   wire n_0_6_13;
   wire n_0_6_14;
   wire n_0_7_0;
   wire n_0_7_1;
   wire n_0_7_2;
   wire n_0_7_3;
   wire n_0_7_4;
   wire n_0_7_5;
   wire n_0_7_6;
   wire n_0_7_10;
   wire n_0_7_11;
   wire n_0_7_12;
   wire n_0_7_13;
   wire n_0_7_14;
   wire n_0_7_7;
   wire n_0_7_9;
   wire n_0_7_8;
   wire n_0_2;
   wire n_0_3;
   wire n_0_5_0;
   wire n_0_5_14;
   wire n_0_5_18;
   wire n_0_5_19;
   wire n_0_5_20;
   wire n_0_5_25;
   wire n_0_5_26;
   wire n_0_5_27;
   wire n_0_5_2;
   wire n_0_5_6;
   wire n_0_5_4;
   wire n_0_5_5;
   wire n_0_5_7;
   wire n_0_5_8;
   wire n_0_5_11;
   wire n_0_5_10;
   wire n_0_5_21;
   wire n_0_5_31;
   wire n_0_5_32;
   wire n_0_5_12;
   wire n_0_5_22;
   wire n_0_5_16;
   wire n_0_5_48;
   wire n_0_5_49;
   wire n_0_5_50;
   wire n_0_5_51;
   wire n_0_5_13;
   wire n_0_5_15;
   wire n_0_5_23;
   wire n_0_5_24;
   wire n_0_5_52;
   wire n_0_5_53;
   wire n_0_5_54;
   wire n_0_5_56;
   wire n_0_5_57;
   wire n_0_5_58;
   wire n_0_5_59;
   wire n_0_5_1;
   wire n_0_5_3;
   wire n_0_5_9;
   wire n_0_5_60;
   wire n_0_5_61;
   wire n_0_5_62;
   wire n_0_5_63;
   wire n_0_5_64;
   wire n_0_1;
   wire n_0_5_28;
   wire n_0_5_29;
   wire n_0_5_67;
   wire n_0_5_30;
   wire n_0_5_71;
   wire n_0_5_72;
   wire n_0_5_73;
   wire n_0_5_33;
   wire n_0_5_34;
   wire n_0_5_35;
   wire n_0_5_36;
   wire n_0_5_37;
   wire n_0_5_38;
   wire n_0_5_39;
   wire n_0_5_40;
   wire n_0_5_41;
   wire n_0_5_42;
   wire n_0_5_43;
   wire n_0_5_45;
   wire n_0_5_65;
   wire n_0_5_66;
   wire n_0_5_68;
   wire n_0_5_69;
   wire n_0_5_70;
   wire n_0_5_74;
   wire n_0_5_75;
   wire n_0_5_76;
   wire n_0_5_77;
   wire n_0_5_78;
   wire n_0_5_79;
   wire n_0_5_80;
   wire n_0_5_83;
   wire n_0_5_85;
   wire n_0_5_86;
   wire n_0_5_87;
   wire n_0_5_89;
   wire n_0_5_17;
   wire n_0_5_44;
   wire n_0_5_46;
   wire n_0_5_47;
   wire n_0_5_55;
   wire n_0_5_81;
   wire n_0_5_82;
   wire n_0_5_84;
   wire n_0_5_88;
   wire [2:0]state;

   INV_X1 i_0_0_0 (.A(ST[1]), .ZN(n_0_0_0));
   INV_X1 i_0_0_1 (.A(ST[2]), .ZN(n_0_0_1));
   INV_X1 i_0_0_2 (.A(ST[3]), .ZN(n_0_0_2));
   INV_X1 i_0_0_3 (.A(n_0_0_3), .ZN(n_0_0));
   NAND2_X1 i_0_0_4 (.A1(n_0_0_4), .A2(n_0_0_6), .ZN(n_0_0_3));
   NAND3_X1 i_0_0_5 (.A1(n_0_0_5), .A2(ST[5]), .A3(ST[4]), .ZN(n_0_0_4));
   NAND3_X1 i_0_0_6 (.A1(n_0_0_1), .A2(n_0_0_0), .A3(n_0_0_2), .ZN(n_0_0_5));
   INV_X1 i_0_0_7 (.A(ST[6]), .ZN(n_0_0_6));
   NOR2_X1 i_0_1_0 (.A1(n_0_1_11), .A2(n_0_1_0), .ZN(alarmbuzz));
   NAND3_X1 i_0_1_1 (.A1(n_0_1_6), .A2(SFA), .A3(n_0_1_1), .ZN(n_0_1_0));
   OAI21_X1 i_0_1_2 (.A(n_0_1_2), .B1(n_0_1_4), .B2(state[2]), .ZN(n_0_1_1));
   NAND3_X1 i_0_1_3 (.A1(n_0_1_10), .A2(n_0_1_9), .A3(n_0_1_3), .ZN(n_0_1_2));
   NAND2_X1 i_0_1_4 (.A1(state[0]), .A2(state[1]), .ZN(n_0_1_3));
   INV_X1 i_0_1_5 (.A(n_0_1_5), .ZN(n_0_1_4));
   NAND3_X1 i_0_1_6 (.A1(SFD), .A2(state[1]), .A3(state[0]), .ZN(n_0_1_5));
   NAND2_X1 i_0_1_7 (.A1(n_0_1_7), .A2(n_0_1_14), .ZN(n_0_1_6));
   OAI211_X1 i_0_1_8 (.A(n_0_1_8), .B(n_0_1_10), .C1(n_0_1_9), .C2(state[0]), 
      .ZN(n_0_1_7));
   NAND2_X1 i_0_1_9 (.A1(SW), .A2(state[1]), .ZN(n_0_1_8));
   INV_X1 i_0_1_10 (.A(SFD), .ZN(n_0_1_9));
   INV_X1 i_0_1_11 (.A(SRD), .ZN(n_0_1_10));
   AOI21_X1 i_0_1_12 (.A(n_0_1_12), .B1(n_0_1_17), .B2(n_0_1_16), .ZN(n_0_1_11));
   OAI21_X1 i_0_1_13 (.A(n_0_1_14), .B1(n_0_1_13), .B2(state[1]), .ZN(n_0_1_12));
   AND2_X1 i_0_1_14 (.A1(n_0_1_15), .A2(state[2]), .ZN(n_0_1_13));
   NAND2_X1 i_0_1_15 (.A1(n_0_1_15), .A2(state[1]), .ZN(n_0_1_14));
   INV_X1 i_0_1_16 (.A(state[0]), .ZN(n_0_1_15));
   INV_X1 i_0_1_17 (.A(n_0_1), .ZN(n_0_1_16));
   INV_X1 i_0_1_18 (.A(n_0_0), .ZN(n_0_1_17));
   XNOR2_X1 i_0_2_0 (.A(state[0]), .B(state[1]), .ZN(n_0_2_0));
   INV_X1 i_0_2_1 (.A(SFA), .ZN(n_0_2_1));
   INV_X1 i_0_2_2 (.A(SRD), .ZN(n_0_2_2));
   INV_X1 i_0_2_3 (.A(SFD), .ZN(n_0_2_3));
   NAND4_X1 i_0_2_4 (.A1(n_0_2_1), .A2(n_0_2_2), .A3(n_0_2_3), .A4(SW), .ZN(
      n_0_2_4));
   NOR2_X1 i_0_2_5 (.A1(n_0_2_0), .A2(n_0_2_4), .ZN(n_0_2_5));
   INV_X1 i_0_2_6 (.A(n_0_3), .ZN(n_0_2_6));
   INV_X1 i_0_2_7 (.A(state[1]), .ZN(n_0_2_7));
   OAI21_X1 i_0_2_8 (.A(n_0_2_7), .B1(SRD), .B2(SFA), .ZN(n_0_2_8));
   NAND2_X1 i_0_2_9 (.A1(n_0_2_8), .A2(SW), .ZN(n_0_2_9));
   NAND2_X1 i_0_2_10 (.A1(n_0_2_7), .A2(SFD), .ZN(n_0_2_10));
   AOI21_X1 i_0_2_11 (.A(state[0]), .B1(n_0_2_10), .B2(n_0_2_1), .ZN(n_0_2_11));
   NOR2_X1 i_0_2_12 (.A1(n_0_2_9), .A2(n_0_2_11), .ZN(n_0_2_12));
   NAND2_X1 i_0_2_13 (.A1(n_0_2_14), .A2(n_0_2_13), .ZN(winbuzz));
   AOI21_X1 i_0_2_14 (.A(n_0_2_5), .B1(n_0_2_12), .B2(n_0_2_6), .ZN(n_0_2_13));
   NAND3_X1 i_0_2_15 (.A1(n_0_2_16), .A2(n_0_2_17), .A3(n_0_2_15), .ZN(n_0_2_14));
   NOR2_X1 i_0_2_16 (.A1(n_0_2_4), .A2(state[0]), .ZN(n_0_2_15));
   INV_X1 i_0_2_17 (.A(n_0_1), .ZN(n_0_2_16));
   INV_X1 i_0_2_18 (.A(n_0_0), .ZN(n_0_2_17));
   INV_X1 i_0_3_0 (.A(state[0]), .ZN(n_0_3_0));
   NAND2_X1 i_0_3_1 (.A1(n_0_3_0), .A2(state[2]), .ZN(n_0_3_1));
   OAI211_X1 i_0_3_2 (.A(n_0_3_1), .B(state[1]), .C1(SW), .C2(state[2]), 
      .ZN(n_0_3_2));
   OAI21_X1 i_0_3_3 (.A(SFD), .B1(state[2]), .B2(state[1]), .ZN(n_0_3_3));
   INV_X1 i_0_3_4 (.A(state[1]), .ZN(n_0_3_4));
   AOI21_X1 i_0_3_5 (.A(n_0_3_5), .B1(n_0_3_12), .B2(n_0_3_11), .ZN(rdoor));
   NAND4_X1 i_0_3_6 (.A1(n_0_3_2), .A2(n_0_3_16), .A3(SRD), .A4(n_0_3_3), 
      .ZN(n_0_3_5));
   NAND2_X1 i_0_3_9 (.A1(SFA), .A2(n_0_3_9), .ZN(n_0_3_6));
   NOR2_X1 i_0_3_10 (.A1(n_0_3_4), .A2(state[2]), .ZN(n_0_3_9));
   INV_X1 i_0_3_11 (.A(state[0]), .ZN(n_0_3_7));
   OAI22_X1 i_0_3_12 (.A1(n_0_3_1), .A2(state[1]), .B1(n_0_3_4), .B2(state[2]), 
      .ZN(n_0_3_11));
   INV_X1 i_0_3_7 (.A(n_0_1), .ZN(n_0_3_8));
   INV_X1 i_0_3_8 (.A(n_0_0), .ZN(n_0_3_10));
   NAND2_X1 i_0_3_13 (.A1(n_0_3_8), .A2(n_0_3_10), .ZN(n_0_3_12));
   INV_X1 i_0_3_14 (.A(n_0_3_7), .ZN(n_0_3_13));
   INV_X1 i_0_3_15 (.A(SFD), .ZN(n_0_3_14));
   AOI21_X1 i_0_3_16 (.A(n_0_3_13), .B1(n_0_3_6), .B2(n_0_3_14), .ZN(n_0_3_15));
   INV_X1 i_0_3_17 (.A(n_0_3_15), .ZN(n_0_3_16));
   INV_X1 i_0_4_1 (.A(state[1]), .ZN(n_0_4_1));
   INV_X1 i_0_4_7 (.A(SW), .ZN(n_0_4_7));
   INV_X1 i_0_4_9 (.A(state[2]), .ZN(n_0_4_9));
   NAND2_X1 i_0_4_0 (.A1(n_0_4_4), .A2(n_0_4_0), .ZN(fdoor));
   NAND2_X1 i_0_4_2 (.A1(SFD), .A2(n_0_4_2), .ZN(n_0_4_0));
   OAI21_X1 i_0_4_3 (.A(n_0_4_3), .B1(n_0_4_13), .B2(state[0]), .ZN(n_0_4_2));
   NAND3_X1 i_0_4_4 (.A1(n_0_4_1), .A2(state[0]), .A3(state[2]), .ZN(n_0_4_3));
   NAND3_X1 i_0_4_5 (.A1(n_0_4_16), .A2(n_0_4_15), .A3(n_0_4_5), .ZN(n_0_4_4));
   AOI21_X1 i_0_4_6 (.A(n_0_4_6), .B1(n_0_4_10), .B2(n_0_4_8), .ZN(n_0_4_5));
   OAI21_X1 i_0_4_8 (.A(SFD), .B1(n_0_4_7), .B2(state[2]), .ZN(n_0_4_6));
   NAND3_X1 i_0_4_10 (.A1(n_0_4_9), .A2(state[0]), .A3(state[1]), .ZN(n_0_4_8));
   OAI21_X1 i_0_4_11 (.A(n_0_4_11), .B1(n_0_4_12), .B2(n_0_4_13), .ZN(n_0_4_10));
   NAND2_X1 i_0_4_12 (.A1(SFA), .A2(n_0_4_9), .ZN(n_0_4_11));
   NOR2_X1 i_0_4_13 (.A1(SRD), .A2(state[2]), .ZN(n_0_4_12));
   XNOR2_X1 i_0_4_14 (.A(n_0_4_14), .B(state[1]), .ZN(n_0_4_13));
   INV_X1 i_0_4_15 (.A(state[2]), .ZN(n_0_4_14));
   INV_X1 i_0_4_16 (.A(n_0_1), .ZN(n_0_4_15));
   INV_X1 i_0_4_17 (.A(n_0_0), .ZN(n_0_4_16));
   NOR2_X1 i_0_6_9 (.A1(SW), .A2(state[2]), .ZN(n_0_6_8));
   OAI21_X1 i_0_6_10 (.A(n_0_6_12), .B1(SFA), .B2(SRD), .ZN(n_0_6_9));
   OAI21_X1 i_0_6_11 (.A(n_0_6_11), .B1(SFA), .B2(n_0_6_12), .ZN(n_0_6_10));
   INV_X1 i_0_6_12 (.A(state[0]), .ZN(n_0_6_11));
   INV_X1 i_0_6_13 (.A(state[1]), .ZN(n_0_6_12));
   INV_X1 i_0_6_0 (.A(n_0_6_0), .ZN(cooler));
   NAND3_X1 i_0_6_1 (.A1(n_0_6_14), .A2(n_0_1), .A3(n_0_6_1), .ZN(n_0_6_0));
   OAI211_X1 i_0_6_2 (.A(n_0_6_2), .B(n_0_6_3), .C1(SW), .C2(n_0_6_4), .ZN(
      n_0_6_1));
   NAND3_X1 i_0_6_3 (.A1(n_0_6_10), .A2(n_0_6_9), .A3(n_0_6_8), .ZN(n_0_6_2));
   NAND3_X1 i_0_6_4 (.A1(n_0_6_11), .A2(n_0_6_12), .A3(state[2]), .ZN(n_0_6_3));
   NAND4_X1 i_0_6_5 (.A1(n_0_6_13), .A2(n_0_6_7), .A3(n_0_6_6), .A4(n_0_6_5), 
      .ZN(n_0_6_4));
   NAND2_X1 i_0_6_6 (.A1(state[0]), .A2(state[1]), .ZN(n_0_6_5));
   INV_X1 i_0_6_7 (.A(SFD), .ZN(n_0_6_6));
   INV_X1 i_0_6_8 (.A(SRD), .ZN(n_0_6_7));
   INV_X1 i_0_6_14 (.A(SFA), .ZN(n_0_6_13));
   INV_X1 i_0_6_15 (.A(n_0_0), .ZN(n_0_6_14));
   INV_X1 i_0_7_0 (.A(n_0_7_0), .ZN(heater));
   NAND2_X1 i_0_7_1 (.A1(n_0_0), .A2(n_0_7_1), .ZN(n_0_7_0));
   OAI21_X1 i_0_7_2 (.A(n_0_7_2), .B1(n_0_7_6), .B2(n_0_7_3), .ZN(n_0_7_1));
   NAND3_X1 i_0_7_3 (.A1(n_0_7_11), .A2(n_0_7_12), .A3(state[2]), .ZN(n_0_7_2));
   OAI21_X1 i_0_7_4 (.A(n_0_7_5), .B1(n_0_7_4), .B2(n_0_7_7), .ZN(n_0_7_3));
   INV_X1 i_0_7_5 (.A(SFA), .ZN(n_0_7_4));
   INV_X1 i_0_7_6 (.A(SW), .ZN(n_0_7_5));
   AOI22_X1 i_0_7_7 (.A1(n_0_7_10), .A2(n_0_7_13), .B1(n_0_7_8), .B2(n_0_7_14), 
      .ZN(n_0_7_6));
   OAI21_X1 i_0_7_8 (.A(n_0_7_12), .B1(SRD), .B2(n_0_7_11), .ZN(n_0_7_10));
   INV_X1 i_0_7_9 (.A(state[0]), .ZN(n_0_7_11));
   INV_X1 i_0_7_10 (.A(state[1]), .ZN(n_0_7_12));
   INV_X1 i_0_7_11 (.A(state[2]), .ZN(n_0_7_13));
   INV_X1 i_0_7_15 (.A(SFD), .ZN(n_0_7_14));
   INV_X1 i_0_7_12 (.A(n_0_7_9), .ZN(n_0_7_7));
   NAND2_X1 i_0_7_13 (.A1(state[0]), .A2(state[1]), .ZN(n_0_7_9));
   AOI21_X1 i_0_7_14 (.A(SRD), .B1(state[0]), .B2(state[1]), .ZN(n_0_7_8));
   INV_X1 i_0_9_0 (.A(Rst), .ZN(n_0_2));
   BUF_X1 rt_shieldBuf__1 (.A(state[2]), .Z(n_0_3));
   NOR2_X1 i_0_5_0 (.A1(SFA), .A2(state[2]), .ZN(n_0_5_0));
   OAI22_X1 i_0_5_1 (.A1(n_0_0), .A2(n_0_5_20), .B1(n_0_5_18), .B2(n_0_5_14), 
      .ZN(display[1]));
   NAND3_X1 i_0_5_2 (.A1(n_0_5_44), .A2(n_0_5_71), .A3(n_0_5_15), .ZN(n_0_5_14));
   AOI21_X1 i_0_5_6 (.A(n_0_5_23), .B1(n_0_5_19), .B2(n_0_5_85), .ZN(n_0_5_18));
   INV_X1 i_0_5_7 (.A(n_0_5_0), .ZN(n_0_5_19));
   AOI21_X1 i_0_5_8 (.A(n_0_5_37), .B1(n_0_1), .B2(n_0_5_43), .ZN(n_0_5_20));
   AOI21_X1 i_0_5_14 (.A(n_0_5_11), .B1(n_0_5_5), .B2(n_0_5_25), .ZN(display[2]));
   NOR2_X1 i_0_5_3 (.A1(n_0_1), .A2(n_0_5_26), .ZN(n_0_5_25));
   AOI21_X1 i_0_5_4 (.A(n_0_5_13), .B1(n_0_5_27), .B2(n_0_5_83), .ZN(n_0_5_26));
   NAND2_X1 i_0_5_10 (.A1(n_0_5_73), .A2(n_0_5_24), .ZN(n_0_5_27));
   NAND2_X1 i_0_5_5 (.A1(SFA), .A2(n_0_5_85), .ZN(n_0_5_2));
   INV_X1 i_0_5_12 (.A(SFA), .ZN(n_0_5_6));
   AOI22_X1 i_0_5_9 (.A1(n_0_5_24), .A2(n_0_5_65), .B1(n_0_5_17), .B2(state[0]), 
      .ZN(n_0_5_4));
   INV_X1 i_0_5_27 (.A(n_0_0), .ZN(n_0_5_5));
   NAND2_X1 i_0_5_29 (.A1(n_0_5_71), .A2(n_0_5_38), .ZN(n_0_5_7));
   NAND2_X1 i_0_5_30 (.A1(n_0_5_4), .A2(n_0_5_38), .ZN(n_0_5_8));
   AOI21_X1 i_0_5_31 (.A(n_0_5_78), .B1(n_0_5_7), .B2(n_0_5_8), .ZN(n_0_5_11));
   INV_X1 i_0_5_11 (.A(n_0_5_65), .ZN(n_0_5_10));
   INV_X1 i_0_5_34 (.A(SRD), .ZN(n_0_5_21));
   INV_X1 i_0_5_35 (.A(SW), .ZN(n_0_5_31));
   NAND2_X1 i_0_5_15 (.A1(SFD), .A2(state[2]), .ZN(n_0_5_32));
   INV_X1 i_0_5_13 (.A(state[1]), .ZN(n_0_5_12));
   INV_X1 i_0_5_18 (.A(SFD), .ZN(n_0_5_22));
   AOI21_X1 i_0_5_21 (.A(n_0_5_84), .B1(n_0_5_22), .B2(n_0_5_89), .ZN(n_0_5_16));
   AOI211_X1 i_0_5_22 (.A(state[2]), .B(n_0_5_12), .C1(n_0_5_2), .C2(SW), 
      .ZN(n_0_5_48));
   NOR2_X1 i_0_5_24 (.A1(n_0_5_31), .A2(SFA), .ZN(n_0_5_49));
   OAI21_X1 i_0_5_25 (.A(n_0_5_32), .B1(n_0_5_49), .B2(SRD), .ZN(n_0_5_50));
   AOI211_X1 i_0_5_26 (.A(n_0_5_16), .B(n_0_5_48), .C1(n_0_5_65), .C2(n_0_5_50), 
      .ZN(n_0_5_51));
   NOR2_X1 i_0_5_28 (.A1(n_0_5_51), .A2(n_0_5_58), .ZN(display[0]));
   BUF_X1 i_0_5_16 (.A(n_0_5_31), .Z(n_0_5_13));
   BUF_X1 i_0_5_19 (.A(n_0_5_32), .Z(n_0_5_15));
   BUF_X1 i_0_5_20 (.A(n_0_5_12), .Z(n_0_5_23));
   BUF_X1 i_0_5_17 (.A(n_0_5_22), .Z(n_0_5_24));
   NAND4_X1 i_0_5_33 (.A1(n_0_5_74), .A2(n_0_5_34), .A3(n_0_5_59), .A4(ST[6]), 
      .ZN(n_0_5_52));
   INV_X1 i_0_5_38 (.A(SRD), .ZN(n_0_5_53));
   INV_X1 i_0_5_37 (.A(n_0_5_23), .ZN(n_0_5_54));
   AOI21_X1 i_0_5_40 (.A(n_0_5_53), .B1(n_0_5_54), .B2(n_0_5_81), .ZN(n_0_5_56));
   OAI21_X1 i_0_5_41 (.A(n_0_5_22), .B1(n_0_5_56), .B2(n_0_5_6), .ZN(n_0_5_57));
   AOI21_X1 i_0_5_44 (.A(n_0_0), .B1(n_0_5_52), .B2(n_0_5_57), .ZN(n_0_5_58));
   NAND3_X1 i_0_5_45 (.A1(n_0_5_1), .A2(n_0_5_3), .A3(n_0_5_9), .ZN(n_0_5_59));
   NOR2_X1 i_0_5_46 (.A1(ST[5]), .A2(ST[3]), .ZN(n_0_5_1));
   NAND3_X1 i_0_5_50 (.A1(ST[1]), .A2(ST[2]), .A3(ST[0]), .ZN(n_0_5_3));
   INV_X1 i_0_5_52 (.A(ST[4]), .ZN(n_0_5_9));
   NOR2_X1 i_0_5_62 (.A1(ST[4]), .A2(ST[5]), .ZN(n_0_5_60));
   NAND3_X1 i_0_5_63 (.A1(ST[1]), .A2(ST[0]), .A3(ST[2]), .ZN(n_0_5_61));
   INV_X1 i_0_5_66 (.A(ST[3]), .ZN(n_0_5_62));
   NAND3_X1 i_0_5_67 (.A1(n_0_5_60), .A2(n_0_5_61), .A3(n_0_5_62), .ZN(n_0_5_63));
   NAND2_X1 i_0_5_68 (.A1(n_0_5_63), .A2(ST[6]), .ZN(n_0_5_64));
   INV_X1 i_0_5_69 (.A(n_0_5_64), .ZN(n_0_1));
   INV_X1 i_0_5_57 (.A(n_0_5_71), .ZN(n_0_5_28));
   INV_X1 i_0_5_72 (.A(SFD), .ZN(n_0_5_29));
   NAND2_X1 i_0_5_23 (.A1(n_0_5_17), .A2(n_0_5_29), .ZN(n_0_5_67));
   INV_X1 i_0_5_32 (.A(n_0_5_67), .ZN(n_0_5_30));
   NAND2_X1 i_0_5_70 (.A1(n_0_5_6), .A2(n_0_5_21), .ZN(n_0_5_71));
   NAND2_X1 i_0_5_71 (.A1(n_0_5_6), .A2(n_0_5_21), .ZN(n_0_5_72));
   INV_X1 i_0_5_77 (.A(n_0_5_72), .ZN(n_0_5_73));
   NOR2_X1 i_0_5_54 (.A1(n_0_5_10), .A2(n_0_5_6), .ZN(n_0_5_33));
   NAND2_X1 i_0_5_58 (.A1(n_0_5_45), .A2(n_0_5_33), .ZN(n_0_5_34));
   NAND2_X1 i_0_5_36 (.A1(n_0_5_30), .A2(n_0_5_13), .ZN(n_0_5_35));
   NAND2_X1 i_0_5_39 (.A1(n_0_5_23), .A2(n_0_5_29), .ZN(n_0_5_36));
   AOI21_X1 i_0_5_43 (.A(n_0_5_28), .B1(n_0_5_35), .B2(n_0_5_36), .ZN(n_0_5_37));
   NAND2_X1 i_0_5_47 (.A1(n_0_5_83), .A2(state[2]), .ZN(n_0_5_38));
   INV_X1 i_0_5_42 (.A(SW), .ZN(n_0_5_39));
   NAND2_X1 i_0_5_48 (.A1(n_0_5_69), .A2(n_0_5_24), .ZN(n_0_5_40));
   NAND2_X1 i_0_5_49 (.A1(n_0_5_87), .A2(n_0_5_46), .ZN(n_0_5_41));
   NAND2_X1 i_0_5_51 (.A1(n_0_5_83), .A2(state[2]), .ZN(n_0_5_42));
   NAND3_X1 i_0_5_53 (.A1(n_0_5_40), .A2(n_0_5_41), .A3(n_0_5_42), .ZN(n_0_5_43));
   NAND2_X1 i_0_5_59 (.A1(n_0_5_47), .A2(state[2]), .ZN(n_0_5_45));
   NAND2_X1 i_0_5_60 (.A1(state[1]), .A2(state[0]), .ZN(n_0_5_65));
   NAND2_X1 i_0_5_74 (.A1(state[0]), .A2(state[1]), .ZN(n_0_5_66));
   NAND2_X1 i_0_5_55 (.A1(n_0_5_39), .A2(n_0_5_66), .ZN(n_0_5_68));
   INV_X1 i_0_5_65 (.A(n_0_5_68), .ZN(n_0_5_69));
   INV_X1 i_0_5_61 (.A(n_0_5_83), .ZN(n_0_5_70));
   OAI21_X1 i_0_5_64 (.A(n_0_5_80), .B1(n_0_5_70), .B2(n_0_5_89), .ZN(n_0_5_74));
   NAND2_X1 i_0_5_56 (.A1(n_0_5_17), .A2(state[1]), .ZN(n_0_5_75));
   INV_X1 i_0_5_90 (.A(n_0_5_75), .ZN(n_0_5_76));
   NAND2_X1 i_0_5_91 (.A1(n_0_5_2), .A2(n_0_5_76), .ZN(n_0_5_77));
   INV_X1 i_0_5_92 (.A(n_0_5_77), .ZN(n_0_5_78));
   NAND2_X1 i_0_5_73 (.A1(n_0_5_81), .A2(n_0_5_12), .ZN(n_0_5_79));
   NAND2_X1 i_0_5_75 (.A1(n_0_5_79), .A2(n_0_5_89), .ZN(n_0_5_80));
   INV_X1 i_0_5_76 (.A(n_0_5_82), .ZN(n_0_5_83));
   INV_X1 i_0_5_94 (.A(state[0]), .ZN(n_0_5_85));
   NAND2_X1 i_0_5_80 (.A1(n_0_5_39), .A2(n_0_5_89), .ZN(n_0_5_86));
   INV_X1 i_0_5_82 (.A(n_0_5_86), .ZN(n_0_5_87));
   INV_X1 i_0_5_78 (.A(state[2]), .ZN(n_0_5_89));
   INV_X1 i_0_5_81 (.A(state[2]), .ZN(n_0_5_17));
   INV_X1 i_0_5_84 (.A(n_0_5_16), .ZN(n_0_5_44));
   NAND2_X1 i_0_5_86 (.A1(n_0_5_81), .A2(n_0_5_12), .ZN(n_0_5_46));
   INV_X1 i_0_5_79 (.A(n_0_5_88), .ZN(n_0_5_47));
   INV_X1 i_0_5_83 (.A(state[0]), .ZN(n_0_5_55));
   INV_X1 i_0_5_85 (.A(state[0]), .ZN(n_0_5_81));
   NAND2_X1 i_0_5_87 (.A1(n_0_5_55), .A2(n_0_5_12), .ZN(n_0_5_82));
   NAND2_X1 i_0_5_88 (.A1(n_0_5_55), .A2(n_0_5_12), .ZN(n_0_5_84));
   NAND2_X1 i_0_5_89 (.A1(n_0_5_55), .A2(n_0_5_12), .ZN(n_0_5_88));
   DFFR_X2 \state_reg[1]  (.D(display[1]), .RN(n_0_2), .CK(clk), .Q(state[1]), 
      .QN());
   DFFR_X2 \state_reg[2]  (.D(display[2]), .RN(n_0_2), .CK(clk), .Q(state[2]), 
      .QN());
   DFFR_X2 \state_reg[0]  (.D(display[0]), .RN(n_0_2), .CK(clk), .Q(state[0]), 
      .QN());
endmodule
